BZh91AY&SY(�$ �߀Py���߰����P9�J�F��$��F(��h��hd 4	*�OHh(�=OSA�  h�h$Q��OP @h    ��b�LFCC �#	 &��M���L�T=@�������SITb,$�$�v���؆���(G�JB
1"�

�a�Ag�A��d�3EI�[����8�SX@�W�K��7� �Ƽ���i{�PZ�D�K
�PЉ�Eg! �	
�4�8�2��E&��T&?��z^��a,�����		0�Y�ƉD���&RDSܶ�5D�t*ı��ţ+'|����k�%aQ�#QQ���G�ьi�������-��-67e�D�Kdg����Hv`��K��6&�Ɍa��0�`�[;hI",aӮ0�����2Q��|XǾ�8���9>�3��b�ͧTSJW���vl�o�>Rk����yaKi�.'�G1�v��C����*��PJ_-,�-NF0,�/!�Li�����h�����s�bw�e���v�'��`;��%�"Sh�s��V�% 1T\7�.0������%<�b���N!�l;$(v�&�Fԉ����
G��2��e��+�B��3׳ZyT,�n��*J��;�Gq��7vby�l��a	�_(�Z L����&�
���
t�/FA��v-�F��x�8"�?eD��R�l�%�L#�r^�L�����"��BN.�U�0�.�,[m�@�B�H-�(&��4!Pu�wԆ��D)�W%d��)4r��2��{���Co�$��m�tg;�*������u!�/�a�[>�#��mhKx���|��ӿ�ݝ�`�,	
�NIBQ��tGl�>�fg�@3�_�}d���I/��]���[��^E�ѝ��lUZLa Hi���I+n���^��*�`$q�+1!,hլ�!T�R��dU[*�j�<`KD��V"��rE8P�(�$